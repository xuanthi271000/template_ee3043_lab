module top (
  // input

  // output

);


endmodule : top
